N-Channel and P-Channel FETs Switch Circuit Transient Response
*
* Including model files
*
*.include NTA4001NT1.LIB
.include NTA4153N.REV0.LIB
.include NTR0202PL.REV0.LIB
*
* Components of the scheme
*
R1 0 1 100k
R2 2 3 100k
* R3 - pull-down resistor to prove an output is floating contact when
* XQ2 is closed
R3 4 0 100k
C1 4 0 1p
XQ1 2 1 0 nta4153n
XQ2 4 2 3 ntr0202plt1
VIN 1 0 pulse (0 3.15 2ms 0ns 0ms 5ms 10ms)
VDD 3 0 pwl (0 0 0ms 0 0ms 3.3v 20ms 3.3v)
*
* Transient analysis for 20ms, step size 0.02ms
*
.tran 0.02ms 20ms
*
* Defining the run-time control functions
*
.control
run
*
* Plotting input and output voltages
*
plot v(1) v(4)
.endc
.end
